//rules of the game:
//1)every row should consist of unique elements
//2)every column should consist of unique elements
//3)every 3x3 subgrid should consist of unique elements
//4)all elements should be in range from 1 to 9

ref:- https://www.edaplayground.com/x/a5D2

class sudoku;
  parameter int M = 3;
  parameter int N = M * M;
  rand bit [7:0] cell[N][N]; //represents every box in the 9x9 grid
  bit [7:0] puzzle[N][N]; //puzzle representing sudoku to be solved
  
  //all elem should be between 1 to 9
  constraint cell_elem_cons {foreach(cell[i,j]){
    cell[i][j] inside {[1:9]};}}
    
  //all row elem in 9x9 grid should be unique
  constraint cell_row_cons {foreach(cell[i,j]){
      foreach(cell[i,k]){
        if(j<k){
          cell[i][j] != cell[i][k];}}}}
          
   //all col elem in 9x9 grid should be unique
   constraint cell_col_cons {foreach(cell[i,j]){
            foreach(cell[k,j]){
              if(i<k){
                cell[i][j] != cell[k][j];}}}}
                
   //all elem in all subgrids (3x3) should be unique
   //i/M == k/M && j/M == l/M tells us that "both cells belong to the same M×M block"
   //The idea for this constraint around integer division to make sure cells across two grids are in same block is borrowed from Keisuke's post. ref:- https://cluelogic.com/2015/02/hidden-gems-of-systemverilog-solving-sudoku/
   constraint subgrid_cons {foreach(cell[i,j]){
                  foreach(cell[k,l]){
                    if((i/M == k/M) && (j/M == l/M) && (i!=k || j!=l)){
                      cell[i][j] != cell[k][l];}}}}
                      
   //The cell should copy over value from the puzzle (if specified)
   //If a cell in the puzzle is zero it is not copied over to the cell. (that is assumed to be solved & generated by the solver)
   constraint puzzle_cell_map_cons {foreach(puzzle[i,j]){
                        if(puzzle[i][j] != 0){
                          cell[i][j] == puzzle[i][j];}}}
endclass
                
                
module tb;
  sudoku s1;
  
  initial begin
    s1=new();
    //The puzzle picked is from wikipedia (ref:- https://en.wikipedia.org/wiki/Sudoku)
    //0 represents element to be generated based on solving constraints by the solver. non-zero elements are just copied over from puzzle grid to cell grid.
    s1.puzzle = '{{5,3,0, 0,7,0, 0,0,0},
                  {6,0,0, 1,9,5, 0,0,0},
                  {0,9,8, 0,0,0, 0,6,0},
                  
                  {8,0,0, 0,6,0, 0,0,3},
                  {4,0,0, 8,0,3, 0,0,1},
                  {7,0,0, 0,2,0, 0,0,6},
                  
                  {0,6,0, 0,0,0, 2,8,0},
                  {0,0,0, 4,1,9, 0,0,5},
                  {0,0,0, 0,8,0, 0,7,9}};
    assert(s1.randomize()) else
      $fatal(0,"randomization error");
    
    //debug disp sudoku solution
    foreach(s1.cell[i]) begin
      $write("%d:",i);
      foreach(s1.cell[,j]) begin
        $write("%d\t",s1.cell[i][j]);
      end
      $display;
    end
  end
endmodule
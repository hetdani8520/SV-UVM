//Problem:-

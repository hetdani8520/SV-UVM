//Signal x should remain high or stable until signal y is asserted. Write a property or assertion.
module x_until_y_assertion;
  bit x, y;
  bit clk;
  
  a1:assert property(@(posedge clk) 
                     1'b1 |-> $stable(x) until y) $display("assertion passed at %tns",$time); else
    $warning("assertion failed at %tns",$time);
    
    
  initial begin
    clk=0;
    forever begin
      #5 clk = ~clk;
    end
  end
    
    //dump waves
  initial begin
  $dumpfile("dump.vcd");
  $dumpvars(1);
  end
    
    initial begin
      x=0;
      y=0;
      repeat(5) @(posedge clk);
      x=0;
      y=1;
      @(posedge clk); //passed at 55ns
      repeat(1) @(posedge clk);
      x=0;
      y=0;
      $finish;
    end
    
endmodule